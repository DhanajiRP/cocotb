module he(a,b);
	input a;
	output reg b;
	always_comb
	begin
                b = a;
	end	
endmodule 
